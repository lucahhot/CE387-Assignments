package edgedetect_uvm_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "edgedetect_uvm_globals.sv"
`include "edgedetect_uvm_sequence.sv"
`include "edgedetect_uvm_monitor.sv"
`include "edgedetect_uvm_driver.sv"
`include "edgedetect_uvm_agent.sv"
`include "edgedetect_uvm_scoreboard.sv"
`include "edgedetect_uvm_config.sv"
`include "edgedetect_uvm_env.sv"
`include "edgedetect_uvm_test.sv"

endpackage
