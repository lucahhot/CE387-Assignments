package cordic_uvm_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "cordic_uvm_globals.sv"
`include "cordic_uvm_sequence.sv"
`include "cordic_uvm_monitor.sv"
`include "cordic_uvm_driver.sv"
`include "cordic_uvm_agent.sv"
`include "cordic_uvm_scoreboard.sv"
`include "cordic_uvm_config.sv"
`include "cordic_uvm_env.sv"
`include "cordic_uvm_test.sv"

endpackage
