package fm_radio_uvm_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "fm_radio_uvm_globals.sv"
`include "fm_radio_uvm_sequence.sv"
`include "fm_radio_uvm_monitor.sv"
`include "fm_radio_uvm_driver.sv"
`include "fm_radio_uvm_agent.sv"
`include "fm_radio_uvm_scoreboard.sv"
`include "fm_radio_uvm_config.sv"
`include "fm_radio_uvm_env.sv"
`include "fm_radio_uvm_test.sv"

endpackage