package udp_reader_uvm_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "udp_reader_uvm_globals.sv"
`include "udp_reader_uvm_sequence.sv"
`include "udp_reader_uvm_monitor.sv"
`include "udp_reader_uvm_driver.sv"
`include "udp_reader_uvm_agent.sv"
`include "udp_reader_uvm_scoreboard.sv"
`include "udp_reader_uvm_config.sv"
`include "udp_reader_uvm_env.sv"
`include "udp_reader_uvm_test.sv"

endpackage
